library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
library UNISIM;
use UNISIM.VComponents.all;
use work.ys_sipm_daq_fpga_type.all;

entity decoder_10b8b is port(
	signal pardat : in std_logic_vector(9 downto 0);
	signal linkok : in std_logic;
	signal clk : in std_logic;
	signal sdin : out std_logic_vector(7 downto 0);
	signal charisk : out std_logic;
	signal dispplus : out std_logic;
	signal dispminus : out std_logic;
	signal notintable : out std_logic
); end decoder_10b8b;

architecture Behavioral of decoder_10b8b is

signal ra : std_logic_vector(13 downto 0);
signal rd : std_logic_vector(15 downto 0);

begin

	ra <= pardat(9 downto 0) & "0000";

	RAMB18E1_decoder_10b8b : RAMB18E1
	generic map (
		INIT_00 => X"0800080008000800080008000800080008000800080008000800080008000800",
		INIT_01 => X"0800080008000800080008000800080008000800080008000800080008000800",
		INIT_02 => X"0800080008000800080008000800080008000800080008000800080008000800",
		INIT_03 => X"0800080008000800080008000800080008000800080008000800080008000800",
		INIT_04 => X"080004EE04ED080004EB08000800080008000800080008000800080008000800",
		INIT_05 => X"080001FE01FD080001FB08000800080001F70800080008000800080008000800",
		INIT_06 => X"0800080008000800080008000800080008000800080008000800080008000800",
		INIT_07 => X"08000800080001FC080008000800080008000800080008000800080008000800",
		INIT_08 => X"0800040E040D0800040B08000800080008000800080008000800080008000800",
		INIT_09 => X"0800001E001D041C001B041A0419080000170416041508000413080008000800",
		INIT_0A => X"080000010002040C0004040A0409080000080406040508000403080008000800",
		INIT_0B => X"080008000800011C0800000F0000040708000010001F04140018041204110800",
		INIT_0C => X"0800006E006D0478006B047F0470080000670460046F0800057C080008000800",
		INIT_0D => X"080008000800007C0800007A0079046808000076007504640073046204610800",
		INIT_0E => X"080008000800006C0800006A00690477080000660065047B0063047D047E0800",
		INIT_0F => X"0800080008000800080008000800080008000800080000740800007200710800",
		INIT_10 => X"0800048E048D0800048B08000800080008000800080008000800080008000800",
		INIT_11 => X"0800009E009D049C009B049A0499080000970496049508000493080008000800",
		INIT_12 => X"080000810082048C0084048A0489080000880486048508000483080008000800",
		INIT_13 => X"080008000800019C0800008F0080048708000090009F04940098049204910800",
		INIT_14 => X"080000AE00AD04B800AB04BF04B0080000A704A004AF0800055C080008000800",
		INIT_15 => X"080002BE02BD00BC02BB00BA00B904A802B700B600B504A400B304A204A10800",
		INIT_16 => X"080002A102A200AC02A400AA00A904B702A800A600A504BB00A304BD04BE0800",
		INIT_17 => X"08000800080003BC080002AF02A000A7080002B002BF00B402B800B200B10800",
		INIT_18 => X"080000CE00CD04D800CB04DF04D0080000C704C004CF0800053C080008000800",
		INIT_19 => X"080002DE02DD00DC02DB00DA00D904C802D700D600D504C400D304C204C10800",
		INIT_1A => X"080002C102C200CC02C400CA00C904D702C800C600C504DB00C304DD04DE0800",
		INIT_1B => X"08000800080003DC080002CF02C000C7080002D002DF00D402D800D200D10800",
		INIT_1C => X"080002EE02ED00F802EB00FF00F0080002E700E000EF08000800080008000800",
		INIT_1D => X"08000800080002FC080002FA02F900E8080002F602F500E402F300E200E10800",
		INIT_1E => X"08000800080002EC080002EA02E900F7080002E602E500FB02E300FD00FE0800",
		INIT_1F => X"0800080008000800080008000800080008000800080008000800080008000800",
		INIT_20 => X"0800080008000800080008000800080008000800080008000800080008000800",
		INIT_21 => X"080000FE00FD04FC00FB04FA04F9080000F704F604F5080004F3080008000800",
		INIT_22 => X"080000E100E204EC00E404EA04E9080000E804E604E5080004E3080008000800",
		INIT_23 => X"0800080008000800080000EF00E004E7080000F000FF04F400F804F204F10800",
		INIT_24 => X"0800002E002D0438002B043F0430080000270420042F080005DC080008000800",
		INIT_25 => X"0800023E023D003C023B003A0039042802370036003504240033042204210800",
		INIT_26 => X"080002210222002C0224002A00290437022800260025043B0023043D043E0800",
		INIT_27 => X"080008000800033C0800022F0220002708000230023F00340238003200310800",
		INIT_28 => X"0800004E004D0458004B045F0450080000470440044F080005BC080008000800",
		INIT_29 => X"0800025E025D005C025B005A0059044802570056005504440053044204410800",
		INIT_2A => X"080002410242004C0244004A00490457024800460045045B0043045D045E0800",
		INIT_2B => X"080008000800035C0800024F0240004708000250025F00540258005200510800",
		INIT_2C => X"0800028E028D0098028B009F0090080002870080008F0800019C080008000800",
		INIT_2D => X"080008000800029C0800029A0299008808000296029500840293008200810800",
		INIT_2E => X"080008000800028C0800028A02890097080002860285009B0283009D009E0800",
		INIT_2F => X"0800080008000800080008000800080008000800080002940800029202910800",
		INIT_30 => X"0800006E006D0800006B08000800080008000800080008000800080008000800",
		INIT_31 => X"0800027E027D007C027B007A0079080002770076007508000073080008000800",
		INIT_32 => X"080002610262006C0264006A0069080002680066006508000063080008000800",
		INIT_33 => X"080008000800037C0800026F0260006708000270027F00740278007200710800",
		INIT_34 => X"0800020E020D0018020B001F0010080002070000000F0800011C080008000800",
		INIT_35 => X"080008000800021C0800021A0219000808000216021500040213000200010800",
		INIT_36 => X"080008000800020C0800020A02090017080002060205001B0203001D001E0800",
		INIT_37 => X"0800080008000800080008000800080008000800080002140800021202110800",
		INIT_38 => X"08000800080008000800080008000800080008000800080001FC080008000800",
		INIT_39 => X"0800080008000800080008000800080008000800080008000800080008000800",
		INIT_3A => X"080008000800080008000800080001F708000800080001FB080001FD01FE0800",
		INIT_3B => X"0800080008000800080008000800080008000800080002F4080002F202F10800",
		INIT_3C => X"0800080008000800080008000800080008000800080008000800080008000800",
		INIT_3D => X"0800080008000800080008000800080008000800080008000800080008000800",
		INIT_3E => X"0800080008000800080008000800080008000800080008000800080008000800",
		INIT_3F => X"0800080008000800080008000800080008000800080008000800080008000800",
		READ_WIDTH_A => 18, 
		READ_WIDTH_B => 18, 
		WRITE_WIDTH_A => 18,
		WRITE_WIDTH_B => 18,
		SIM_DEVICE => "7SERIES"
	)
	port map (
		DOADO => rd,
		DOPADOP => open,
		DOBDO => open,
		DOPBDOP => open,
		ADDRARDADDR => ra, 
		CLKARDCLK => clk,
		ENARDEN => linkok,
		REGCEAREGCE => '1',
		RSTRAMARSTRAM => '0',
		RSTREGARSTREG => '0',
		WEA => "00",
		DIADI => "1111111111111111",
		DIPADIP => "11",
		ADDRBWRADDR => "11111111111111",
		CLKBWRCLK => clk,
		ENBWREN => '0',
		REGCEB => '1',
		RSTRAMB => '0',
		RSTREGB => '0',
		WEBWE => "0000",
		DIBDI => "1111111111111111",
		DIPBDIP => "11"
	);

	sdin <= rd(7 downto 0);
	charisk <= rd(8);
	dispplus <= rd(9);
	dispminus <= rd(10);
	notintable <= rd(11);

end Behavioral;

